
`include "time_sleuth/defines.v"

import my_types::*;

module resolution(
    input clock,
    input VideoMode videoMode,
    input [3:0] addr,
    output [`RESLINE_SIZE-1:0] q
);

    reg [`RESLINE_SIZE-1:0] q_reg;

    always @(posedge clock) begin
        case (addr)
            00: q_reg <= 0;
            01: q_reg <= 0;
            02: q_reg <= { 96'b111111100001000000000000000000000000000000111100000100000000000000000000000100000100000000000000, (videoMode.id[3] ? 32'b00000000000010000011110000111100 : (videoMode.id[2] ? 32'b00000000011111100011110000111100 : 32'b00011000001111000011110000111100)), (videoMode.id[0] ? 8'b00010000 : 8'b00000000 ) };
            03: q_reg <= { 96'b000100000000000000000000000000000000000001000010000100000000000000000000000100000100000000000000, (videoMode.id[3] ? 32'b00000000000010000100001001000010 : (videoMode.id[2] ? 32'b00000000000000100100001001000010 : 32'b00101000010000100100001001000010)), (videoMode.id[0] ? 8'b00000000 : 8'b00000000 ) };
            04: q_reg <= { 96'b000100000000000000000000000000000000000001000000000100000000000000000000000100000100000000000000, (videoMode.id[3] ? 32'b00000000000110000100001001000010 : (videoMode.id[2] ? 32'b00000000000000100000001001000010 : 32'b00001000010000100100001001000010)), (videoMode.id[0] ? 8'b00000000 : 8'b00000000 ) };
            05: q_reg <= { 96'b000100000011000001101000001110000000000001000000000100000011100001000100001110000111100000000000, (videoMode.id[3] ? 32'b00000000000110000100001001000110 : (videoMode.id[2] ? 32'b00000000000001000000001001000110 : 32'b00001000010001100100001001000110)), (videoMode.id[0] ? 8'b00110000 : 8'b01111000 ) };
            06: q_reg <= { 96'b000100000001000001010100010001000000000000111100000100000100010001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000001010000011110001001010 : (videoMode.id[2] ? 32'b00000000000001000000001001001010 : 32'b00001000010010100011110001001010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            07: q_reg <= { 96'b000100000001000001010100010001000000000000000010000100000100010001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000001010000100001001010010 : (videoMode.id[2] ? 32'b00000000000010000000001001010010 : 32'b00001000010100100100001001010010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            08: q_reg <= { 96'b000100000001000001010100011110000000000000000010000100000111100001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000010010000100001001100010 : (videoMode.id[2] ? 32'b00000000000010000011110001100010 : 32'b00001000011000100100001001100010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            09: q_reg <= { 96'b000100000001000001010100010000000000000000000010000100000100000001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000010010000100001001000010 : (videoMode.id[2] ? 32'b00000000000100000100000001000010 : 32'b00001000010000100100001001000010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            10: q_reg <= { 96'b000100000001000001010100010000000000000000000010000100000100000001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000011111100100001001000010 : (videoMode.id[2] ? 32'b00000000000100000100000001000010 : 32'b00001000010000100100001001000010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            11: q_reg <= { 96'b000100000001000001010100010000000000000001000010000100000100000001000100000100000100010000000000, (videoMode.id[3] ? 32'b00000000000010000100001001000010 : (videoMode.id[2] ? 32'b00000000000100000100000001000010 : 32'b00001000010000100100001001000010)), (videoMode.id[0] ? 8'b00010000 : 8'b01000100 ) };
            12: q_reg <= { 96'b000100000011100001010100001111000000000000111100000011000011110000111000000011000100010000000000, (videoMode.id[3] ? 32'b00000000000010000011110000111100 : (videoMode.id[2] ? 32'b00000000000100000111111000111100 : 32'b00111110001111000011110000111100)), (videoMode.id[0] ? 8'b00111000 : 8'b01111000 ) };
            13: q_reg <= { 128'b0, (videoMode.id[0] ? 8'b00000000 : 8'b01000000 ) };
            14: q_reg <= { 128'b0, (videoMode.id[0] ? 8'b00000000 : 8'b01000000 ) };
            15: q_reg <= { 128'b0, (videoMode.id[0] ? 8'b00000000 : 8'b01000000 ) };
        endcase
    end

    assign q = q_reg;

endmodule 


